`timescale 1ns / 1ps
module seven_segment(
    );


endmodule